module ubus_tb_top;
    import uvm_pkg::*;

    initial begin
        run_test();
    end
endmodule : ubus_tb_top