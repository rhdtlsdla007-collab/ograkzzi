package jk_ubus_common_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"


  
endpackage : jk_ubus_common_pkg

