class test;

endclass