package router_stimulus_pkg;

import uvm_pkg::*;

`include "packet.sv"

 
 
 
`include "packet_sequence.sv"




 
 
 
`include "packet_da_3.sv"






endpackage
