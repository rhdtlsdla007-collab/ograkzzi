package jk_ubus_common_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"


  `include "../slave/jk_ubus_slave_transfer.sv"
endpackage : jk_ubus_common_pkg

