class jk_ubus_test extends uvm_test;
    `uvm_component_utils(jk_ubus_test)
    jk_ubus_env env;

    function new(string name, uvm_component parent);
    super.new(name, parent);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
    endfunction: new

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        env = jk_ubus_env::type_id::create("env", this);
        uvm_config_db#(uvm_object_wrapper)::set(this, "env.master_agent.sqr.run_phase", "default_sequence", jk_ubus_master_sequence::type_id::get());
        uvm_config_db#(uvm_object_wrapper)::set(this, "env.slave_agent.sequencer.run_phase", "default_sequence", jk_ubus_slave_sequence::type_id::get());
    endfunction

    function void end_of_elaboration_phase(uvm_phase phase);
        uvm_top.print_topology();
    endfunction

    task run_phase(uvm_phase phase);
        phase.raise_objection(this);
            #1000ns;
        phase.drop_objection(this);
    endtask
endclass : jk_ubus_test

/////////////////////////

class jk_ubus_virtual_sequence_test extends uvm_test;
 `uvm_component_utils(jk_ubus_virtual_sequence_test)

 jk_ubus_env env;
 jk_ubus_virtual_sequence virtual_sequence;

 function new(string name = "jk_ubus_virtual_sequence_test", uvm_component parent = null);
	super.new(name, parent);
 endfunction

 function void build_phase(uvm_phase phase);
	super.build_phase(phase);
	env = jk_ubus_env::type_id::create("env", this);
 endfunction

 function void end_of_elaboration_phase(uvm_phase phase);
	uvm_top.print_topology();
 endfunction

 task run_phase(uvm_phase phase);
	phase.raise_objection(this);
	virtual_sequence = jk_ubus_virtual_sequence::type_id::create("virtual_sequence");
	virtual_sequence.start(env.virtual_sequencer);
	phase.drop_objection(this);
 endtask

endclass : jk_ubus_virtual_sequence_test

