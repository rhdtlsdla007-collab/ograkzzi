class jk_ubus_virtual_sequencer extends uvm_sequencer;
 `uvm_component_utils(jk_ubus_virtual_sequencer)

 function new(string name = "jk_ubus_virtual_sequencer", uvm_componenet parent=null);
	super.new(name, parent);
 endfunction

endclass

